// Code your design here
/*what is Fibonacci series/sequence.
  The Fibonacci series is a series of non-negative integers where an element is the addition of the two previous elements of the series.
The first two elements are pre-defined: 
  						f[0] = 0 and f[1] = 1.
All subsequent elements for (n >= 2) are f[n] = f[n-1] + f[n-2].
Thus, the first few elements of the Fibonacci series are:
  							0, 1, 1, 2, 3, 5, 8, 13, 21, 34, 55…*/