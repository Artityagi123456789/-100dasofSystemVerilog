module tb;
int array;
initial begin
	array = 8'b0101010101;
	for(i=0;i<size(array);i++)begin
	$display("value of arr_data[i]);

	end
end
endmodule
